module IC90_TB;

    // Inputs
    reg cka;
    reg ckb;
    reg r0_1;
    reg r0_2;
    reg r9_1;
    reg r9_2;

    // Outputs
    wire [3:0] q;

    // Instantiate the Unit Under Test (UUT)
    IC90 uut (
        .cka(cka),
        .ckb(ckb),
        .r0_1(r0_1),
        .r0_2(r0_2),
        .r9_1(r9_1),
        .r9_2(r9_2),
        .q(q)
    );

    // Clock generation for cka (divide-by-2 section)
    initial begin
        cka = 0;
        forever #5 cka = ~cka; // Toggle cka every 5 ns
    end

    // Clock generation for ckb (divide-by-5 section)
    initial begin
        ckb = 0;
        forever #10 ckb = ~ckb; // Toggle ckb every 10 ns
    end

    // Test sequence
    initial begin
        // Initialize inputs
        r0_1 = 1;
        r0_2 = 1;
        r9_1 = 1;
        r9_2 = 1;

        // Apply asynchronous reset to start from 0
        #10 r0_1 = 0; r0_2 = 0; // Apply reset
        #10 r0_1 = 1; r0_2 = 1; // Release reset

        // Wait to observe the counter increment
        #200;

        // Test reset when counter reaches 9
        #10 r9_1 = 0; r9_2 = 0; // Apply reset
        #10 r9_1 = 1; r9_2 = 1; // Release reset

        // Wait to observe the counter reset and start over
        #200;

        // Finish simulation
        $finish;
    end

    // Monitor outputs
    initial begin
        $monitor("Time = %0dns, cka = %b, ckb = %b, r0_1 = %b, r0_2 = %b, r9_1 = %b, r9_2 = %b, q = %b", 
                 $time, cka, ckb, r0_1, r0_2, r9_1, r9_2, q);
    end

endmodule
