module IC76(
    input clk,
    input reset,
    input set,
    input j, k,
    output reg q,
    output q_inverted
);

    // Assign the inverted output
    assign q_inverted = ~q;

    // Always block triggered on the negative edge of clk
    always @(negedge clk) begin
        if (reset) begin
            q <= 1'b0; // Asynchronous reset to 0
        end else if (set) begin
            q <= 1'b1; // Asynchronous set to 1
        end else begin
            case ({j, k}) // Concatenate j and k to form a 2-bit value
                2'b00: q <= q;      // No change
                2'b01: q <= 1'b0;   // Reset
                2'b10: q <= 1'b1;   // Set
                2'b11: q <= ~q;     // Toggle
            endcase
        end
    end
endmodule
